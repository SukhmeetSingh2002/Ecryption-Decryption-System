module bit_rand_11 (rand_11);
    output [10:0]rand_11;
    reg [10:0]rand_11;
    
endmodule