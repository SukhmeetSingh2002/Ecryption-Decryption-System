module bit_rand_9 RAND1(rand_9);
    output [8:0]rand_6;
    reg [8:0]rand_6;
    
endmodule