module bit_rand_6 RAND1(rand_6);
    output [5:0]rand_6;
    reg [5:0]rand_6;
    
endmodule