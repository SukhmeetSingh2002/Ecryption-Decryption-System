module 6_bit_rand RAND1(Clk,6_rand);
    input Clk;
    output [5:0]6_rand;
    reg [5:0]6_rand;
endmodule